package router_pkg;

	import uvm_pkg::*;

	`include "uvm_macros.svh"
	
	`include "source_xtn.sv"
	`include "source_config.sv"
	`include "destination_config.sv"
	`include "env_config.sv"
	`include "source_driver.sv"
	`include "source_monitor.sv"
	`include "source_sequencer.sv"
	`include "source.sv"
	`include "router_source_top.sv"
	`include "source_sequence.sv"
	
	`include "destination_xtn.sv"
	`include "destination_monitor.sv"
	`include "destination_sequencer.sv"
	`include "destination_sequence.sv"		
	`include "destination_driver.sv"
	`include "destination.sv"
	`include "router_destination_top.sv"
	
	`include "router_scoreboard.sv"
	`include "env.sv"

	`include "test.sv"




endpackage
